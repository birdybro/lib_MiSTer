    INIT_00 => x"FBFC1BFD18FA18FA18FA18FA18FA4FFC53FC5EFCABFC65FCA9FC80FC7CF838F8",
    INIT_01 => x"C6C0F08E10B9FE8EC0F0CE100CFD04FDFBFCFAFCEBFCDCFCD2FCBFFC3AFD04FD",
    INIT_02 => x"A7D0866AAFDD8C30FB265AE26F0CC68E0117D0F0BF00E08EF9265AA0A780A610",
    INIT_03 => x"17E5FE8EE20317C9FE8EA504178704174F0417D8F0B70386D7F0B70386431FE4",
    INIT_04 => x"A302170E0417408B981F1504175E86092C2081891FF1270D817F84FB0317CD03",
    INIT_05 => x"1F2D29450217C22094ADC620AA0317E7FE8EF526B9FE8C02300F2780E17AFE8E",
    INIT_06 => x"E127088111283802176C0217650317A4A6740217650317211F880317EDFE8E12",
    INIT_07 => x"31C2202131B003173F864D02170827A4A1A4A7390F260D8117275E81DD271881",
    INIT_08 => x"1000C3101F390124E1AC20340629E6011705201F30C0F08E321FC00217BE203F",
    INIT_09 => x"E4AE110317EDFE8E103439623203273403170527E4AC011FF0C4201F0634F0C4",
    INIT_0a => x"0425208180A610C6E1AEEB0117F5265AF30117EC021780A610C6FB0117EE0217",
    INIT_0b => x"17072653810503175F3B341F390128FD0117BC20EE265A4203172E8602237E81",
    INIT_0c => x"1F031707265381E702175F39D7F0F7E72001C88E031707265681F22002C83D03",
    INIT_0d => x"8E10341A24C0F08C1E294C011739D8F0F7E72001C84F031707264B81F22002C8",
    INIT_0e => x"10CC02163F866901173984A73F86A4AFA0A709273F8184A60F271035558DFFFF",
    INIT_0f => x"AE7DFE16AC0117068D4AAF0427268D1F304AAE431F39FB265A188D08C6D9F08E",

    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000",

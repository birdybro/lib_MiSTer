    INIT_00 => x"A608C6D9F08E1039A0A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0F08C21",
    INIT_01 => x"273981670217F92653816E0217D2F07F528D1186393D3139F7265A0427A1ACA0",
    INIT_02 => x"170434E46AE46AE4EBE0EBE0E610342129B3001726290234CA0017F12631813C",
    INIT_03 => x"D2F073058D3F86B327FFC102355FEB2080A70527E46AE0EB02340C290435B000",
    INIT_04 => x"062762A3E4EC1102171286E4AF0130462562AC4A2930346F8DE26F2602161386",
    INIT_05 => x"63EB62EB75011762AE820117981F03CB9F01172EFF8E64E720C6022320008310",
    INIT_06 => x"188D3965326A8D1486C326E4AC62AF680117981F53F526646A72011780A684EB",
    INIT_07 => x"2D86121F4229088D391035F726E4AC1080A7A0A60929188D5D8D3E8610341529",
    INIT_08 => x"1E29078D891F484848482829118D903561A710343229088D011F38290E8D438D",
    INIT_09 => x"021A393780032246810725418139308003223981122530817C011739E0AB0434",
    INIT_0a => x"3941A70229B78DEA8D8300173944AF0229B38DF68D8500176301162086008D39",
    INIT_0b => x"AF0229858DC88D7C8D394AAF0229908DD38D7E8D3943A70229AB8DDE8D800017",
    INIT_0c => x"FF17A58D748D3942A702297DFF17B18D778D3946AF022979FF17BD8D7A8D3948",
    INIT_0d => x"358D910017EDFE8E348D2D8D268D1E8D168DA10017EDFE8E39C4A7808A042971",
    INIT_0e => x"A67F8D15FF8E572044AE88001709FF8E6120311F920017F1FE8E4A20438D3C8D",
    INIT_0f => x"FF8E332048AE648DFDFE8E3C204AAE6D8DF7FE8E4D2043A6768D0FFF8E562041",

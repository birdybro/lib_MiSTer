    INIT_00 => x"50814CD3F0FC3903E702A7D3F0FDD4F0F64F39D6F07FF726508102A74C84E720",
    INIT_01 => x"A702E7D3F0F72086D3F0F604E75F012519C15C04E6E78D5AEA2619C15C4FF026",
    INIT_02 => x"39D6F0F702E7D3F0F75FE4205F03E7D4F0F7082719C15CD4F0F6F42650C15C84",
    INIT_03 => x"8EFB0254FB01E62073FE178FFE17EE20CAFE176FFE17F6276AFE170D2698FE17",
    INIT_04 => x"F9496EF9470FF945B3F94260FE4182FB1948FB1877FB156CFB1060FB049AFB03",
    INIT_05 => x"F976F976F976F9DEFA5ADFF95803F953A8FB5285FA5077F94FBAF84D2CFA4C95",
    INIT_06 => x"0D0420302E31562053394755422D4B0000000A0D000000FFFFFFFFEBF976F976",
    INIT_07 => x"552020043D43502020043D5053202004202D20043F54414857043E040000000A",
    INIT_08 => x"20043D422020043D412020043D50442020043D58492020043D59492020043D50",
    INIT_09 => x"00000000000000000000000000000004315343565A4E4948464504203A434320",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"9F6EC6F09F6EC4F09F6EC0F09F6E000000000000000000000000000000000000",
    INIT_0e => x"0822CEF0BC8B300F27FFFF8CCCF0BE49584F4AAF80E64AAE431FCAF09F6EC8F0",
    INIT_0f => x"34F834F8C2FFBEFFBAFFB6FFC6FFB2FFC2F09F6E42EE1F37F16E44AEC4EC1034",

    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_11 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_12 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_13 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_14 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_15 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_16 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_17 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_21 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_22 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_23 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_24 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_25 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_26 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_27 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_28 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_29 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_2f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_30 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_31 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_32 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"0000000000000000000000000000000000000000000000000000000000000000",

    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000E4CC7E",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"00000000000000000000000000000000005458540050555452415453000000FF",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_10 => x"CDBFFBD3BEF1D39FAD06CABFA10089302BCCBEFDD3B73986A0C039ACCABD0620",
    INIT_11 => x"2684E11284E784A6B9C6A0008E4FCDBFF7D3BE13CDBF10CDBFF9D3BE0DCDBF0A",
    INIT_12 => x"BD81CEBDDCCA8E16CCBF03CD8E2BCCBF5FFF8930EC2606CABC0004893084A70B",
    INIT_13 => x"CCBF80C08E67CD7E00D2BD01A6082706D4BD84A7018640C88EB5CEBD9E8DB5CE",
    INIT_14 => x"80C08EF4D1BD40C88EE7260D8180A714CCBED7D27E3034052706D4BD40C88E14",
    INIT_15 => x"EC250D8D0ECCB7F325148D2BCEBD81CEBDECCA8E2ED37E43CCBF67CD8E14CCBF",
    INIT_16 => x"3930383639011A39FE1C03275D1CCCB60B2575D1BD3910CCB7E525068D0FCCB7",
    INIT_17 => x"000004203F2959592C44442C4D4D2820455441440431302E33562058454C4620",
    INIT_18 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_19 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_1f => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_20 => x"0000000000000000000000000000000000000001001BFF0000400400193A1808",
    INIT_21 => x"00000000000000000000000000000000010000FFBF0000000000000000000000",
    INIT_22 => x"274E4143043F54414857043F3F3F042B2B2B0000000060000000000000000000",
    INIT_23 => x"20524F525245204B53494404444E554F4620544F4E04524546534E4152542054",
    INIT_24 => x"004BD3004E4F4D0FD20054454704594441455220544F4E205345564952440423",
    INIT_25 => x"0000000000000000000000000000000000000000000000000A006400E8031027",
    INIT_26 => x"000000000070D37E00000000000000000000000000000000000000000070D37E",
    INIT_27 => x"0000000000000001000000000000000000000000000000000070D37E00000000",
    INIT_28 => x"CE7E2BCE7E41CF7EFBCE7E12CD7E0FCD7E0CCD7E09CD7EB1CD7E67CD7E57CD7E",
    INIT_29 => x"7ED4CF7E86CF7E49D37EEBD07EA2D17E36D07EEACD7E0ED07EB5CE7EEDCF7E81",
    INIT_2a => x"D4BD11CC7F7FC0CE1005CE7E05CE7E4ECD7E29D37E75D17ED0CF7E2FD17E7FD2",
    INIT_2b => x"9FAFE7D3BEE9D39FAF00C78E16CCBF03CD8E18DEBD7FC0CE10FDD3BD28CC7F00",
    INIT_2c => x"28CC7D142015CC7C052602CCB111CCB65A8D4CCC7F34CC7F31CCBFF8CC8EEBD3",
    INIT_2d => x"D0BD0DCC7C40C88EE5270D81D4D0BD7A8D81CEBD4ECC8EB22603D4BD97052610",
    INIT_2e => x"CCB7158656CC8E2ED2BD01986E0326358D072712CCBE09273E8D93CC8E162536",
    INIT_2f => x"7F21CC7F22CC7F23CC7F0ACDBF0DCDBE10CDBF13CDBE67CD7E11CC7F81CEBD20",
    INIT_30 => x"806D0C27A46DF026846D082680A1208002235F81A0A644C88E103924CC7F26CC",
    INIT_31 => x"0D811F2700CCB11D2701CCB1FBCEBD14CCBF80C08E39FB1CDE26846D0230FC26",
    INIT_32 => x"80C08CCE20268D52CC8E39DC260D8180A7E227FFC08CE7231F8132270A810D27",
    INIT_33 => x"20208641CFBD0D86B92066CFBD07CCB666CFBD20860826088107CCB61F30F427",
    INIT_34 => x"CC7F5C26121381E5D39FAD65274ECDBDF320013041CFBD6F27048184A6328DC9",
    INIT_35 => x"2703CCB6D48D272621CC7D16CC9F6E11CC7FF32603815027121181E5D39FAD1A",
    INIT_36 => x"CC7C0435FB265A088D052708CCF60434CE8D022709CC7D1ACC7F18221ACCB120",
    INIT_37 => x"1A2623CC7D39FE1C0435FA265A4E8D4F062705CCF60434588D0A865C8D0D861A",
    INIT_38 => x"1ACC7F0CCDBD032009CDBD0820538D0C2724CC7D11272FCC7D1A8D102726CC7D",
    INIT_39 => x"CD7E7FD2BD24CC7F3947CCBE042606D4BD24CCBE47CCBF062026CCBE47CCBF39",
    INIT_3a => x"CEBD062429CCB10B2704CCB6023429CC7C172029CC7F05221F81202621CC7D03",
    INIT_3b => x"03200FCDBD082626CC7D0D20B58D042724CC7D132622CC7D0234023529CC7CB5",
    INIT_3c => x"1FF7264DCC7A02300B8DA0CC8E84EC4DCCB704861DCCF74ACC7F39023512CDBD",
    INIT_3d => x"CC7D0B264ACC7D10264BCCB60234F4204BCC7C84A3072584A3104BCC7F3D2098",
    INIT_3e => x"44444444042084A6048D84A60130028D8235128D4ACC7C0520238D20860B271D",
    INIT_3f => x"2561810E235A810C254181162339811425308141CF7E078B02233981308B0F84",

    INIT_00 => x"063428F6F629F6B6063426F6F627F6B6063424F6F625F6B606342EF6F62FF6B6",
    INIT_01 => x"1022F6F723F6B7401F3B0234508A2DF6B602342BF6B602342AF6B602342CF6B6",
    INIT_02 => x"A4A6021F01E602A6043420275454C0A7008631F6CED1FD7E21F6B7008620F6CE",
    INIT_03 => x"A6021F84E601A69CFE7EE02631F6F1043031F67CC0A70C260435A4E1A4E703E6",
    INIT_04 => x"40B4FEBD002031F6B7018632F6B792FE7E4FA4A702A6021F84E601A692FE7EA4",
    INIT_05 => x"5A80AB008602CB01E630F68EF1FC7EF8265A7CFCBD80A603CB01E630F68E84A7",
    INIT_06 => x"26508502352BF6B7846E04F0BE0586846E02F0BE0686846E00F0BE078639FB26",
    INIT_07 => x"6E0CF0BE0286846E08F0BE0386846E06F0BE04860234508A04342BF6F67C3409",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000ACFC7E018684",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0f => x"00FCFAFE01FFF3FED8FED1FECAFEC3FE00000000000000000000000000000000",

    INIT_00 => x"A0E8E0EB023464E3201F62AE10F125E4AC10A0A7E0AB043464E3201FE8031777",
    INIT_01 => x"3903175003174701171035880317A1FE8E10344C03173F3085031783FE8E3C27",
    INIT_02 => x"AC101A268303173E0317A6FE8E981F6C03178FFE8E2E031764AE77031787FE8E",
    INIT_03 => x"1E29B102173966328C26646C9026656C62AE100B267403178603172B86B325E4",
    INIT_04 => x"173984A73F86A4AFA0A709273F8184A60F271035558DFFFF8E10341A24C0DF8C",
    INIT_05 => x"8D4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF8E104703163F864A03",
    INIT_06 => x"A0A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C21AE9AFD16E4FD1706",
    INIT_07 => x"F0B714F0B7FF8624F0B7DE86393D3139F7265A0427A1ACA0A608C6E3DF8E1039",
    INIT_08 => x"B68A001720F0B70986FB2B20F0B697001720F0B7D88610F07D16F0B715F0B710",
    INIT_09 => x"F0BFFFFE8E00F0FD5343101F40F0B7108A528D00C08ECA261085F926018520F0",
    INIT_0a => x"0A2A10F07D5F04345F528D20F0B78C8622F0B7018614F0B7FE8610F0B7FF8602",
    INIT_0b => x"341F4AAF00C08E24F0F7DEC63901271C8520F0B604358A20F0265A0435F8265A",
    INIT_0c => x"0F8462A65858585853A6E6E4E754545454A6E6D0DF8E104444444462A636343B",
    INIT_0d => x"013000008E03C614E07F18E07D390435FD265A20C6043439363562E762EA62A7",
    INIT_0e => x"B78C86298D1AE0B70186F92601C518E0F6378D18E0B70F86F6265AF92600008C",
    INIT_0f => x"C08E3901272CC5F02601C518E0F680A71BE0B6052702C5092000C08E228D18E0",

    INIT_00 => x"2650C15C84A702E7FBDFF72086FBDFF604E75F012519C15C04E6E78D5AEA2619",
    INIT_01 => x"FB0274FB0139FEDFF702E7FBDFF75FE4205F03E7FCDFF7082719C15CFCDFF6F4",
    INIT_02 => x"505EFA4CA5F847FDF8455CF94248FB1953FB183DFB1531FB105EFB047FFB0369",
    INIT_03 => x"94F9A7F8A7F8A7F8A7F894F992FC55D5F94488F958F1F853EDFB52A8F84DBCFA",
    INIT_04 => x"20204147504620524F4620322E312047554239305359530000000A0DFFFFFFFF",
    INIT_05 => x"43502020043D5053202004202D20043F54414857043E040000000A0D4B04202D",
    INIT_06 => x"20043D412020043D50442020043D58492020043D59492020043D53552020043D",
    INIT_07 => x"0000000000000000000004315343565A4E4948464504203A43432020043D4220",
    INIT_08 => x"300B2784AC1084AF1084EEAA558E10A0D08E84A7F086FB264A80A70F86F0FF8E",
    INIT_09 => x"2DA7D0DF8E10C0DFCE10FDFFB74444444443101F84EFD620ED26A0F08C00F089",
    INIT_0a => x"1084AF10AA558E1084EE2227A0F08C00F08930FB2A4AA66F0C862FA7F0862E6F",
    INIT_0b => x"2EA7D0DF8E10F186D520A5A70F88891F44444444101FD0DF8E1084EFE92684AC",
    INIT_0c => x"8EF32D0C814C80E7A66F0427A6E6211F4F2CE7A66F1420F92A4A0526A6E60C86",
    INIT_0d => x"9F6EC6DF9F6EC4DF9F6EC0DF9F6E62F816E2DFF753F9265A80A7A0A610C6F0FF",
    INIT_0e => x"0822CEDFBC8B300F27FFFF8CCCDFBE49584F4AAF80E64AAE431FCADF9F6EC8DF",
    INIT_0f => x"00FFB2FFC2FFBEFFBAFFB6FFC6FFB2FFC2DF9F6E42EE1F37F16E44AEC4EC1034",

    INIT_00 => x"3FF13FF13FF141F119F152F052F052F03FF13FF13FF13FF13FF141F119F1BDF7",
    INIT_01 => x"7AF152F052F052F052F052F052F052F052F052F052F052F052F052F03FF13FF1",
    INIT_02 => x"6E34DE9F6E32DE9F6E39FE1C5D5F52F052F052F04EF24EF24EF24EF249F2E9F1",
    INIT_03 => x"0FC630350826FF8185A62ADE8E1EDEF703E6303438DE9F6E390127078D36DE9F",
    INIT_04 => x"6E3ADE9F6E3035F9265AA0A780A614C632DE8E108B3002F08E3D14C639011A5D",
    INIT_05 => x"6E39EA2604814C1EDEB640DE9FAD0425BC8D1BDE8E1EDEB74F3EDE9F6E3CDE9F",
    INIT_06 => x"F084C5AB1FDEB62EDECEC5E61EDEF62ADECE501A22DEB7A81F44DE9F6E42DE9F",
    INIT_07 => x"B70F88008639031F5F008B0F841FDEB6F0FFB7E0AB0F840F88018020DEB6E2A7",
    INIT_08 => x"FF17EAFF17703439011A5D40C639041AFE1C20DEF71FDEB7398A1F22DEB6F0FF",
    INIT_09 => x"5FF0355FF9265A80A7A0A65F46DE8E10CBFF17F9265AA0A7C0A65F46DE8E10A6",
    INIT_0a => x"80A65F46DE8E10BAFF16032700C1072701C1C5E61EDEF62ADECEC2FF17703439",
    INIT_0b => x"DE7F02340434F0355F84FF17F9265AC0A7A0A65F46DE8E105FFF17F9265AA0A7",
    INIT_0c => x"2485F2BD02353D2485F2BD0235442485F2BD1EDEB64C2485F2BD738622DE7F21",
    INIT_0d => x"F2BD02341B2467F2BDEB265A21DE7C032422DEB722DEBB80A7302467F2BD5F36",
    INIT_0e => x"85F2BD1586092010C60D205F032485F2BD06860E2621DEB3100235891F142467",
    INIT_0f => x"85F2BD1EDEB6DD2485F2BD728622DE7F21DE7F02340434395D21DEF709C6F524",
    INIT_10 => x"032422DEB722DEBBBF2485F2BD80A65FC72485F2BD0235CE2485F2BD0235D524",
    INIT_11 => x"5F032606819C2467F2BDA12485F2BD22DEB6A92485F2BD21DEB6EB265A21DE7C",
    INIT_12 => x"205F03260681072467F2BD0C2485F2BD5186395D21DEF6395D21DEF70AC60220",
    INIT_13 => x"B035EE261F30F6263F310A254700E0B6E2048E10E8038E3034395D011A10C604",
    INIT_14 => x"35ED261F30F5263F310C25474700E0B6E2048E10E8038E02343034B03501E0B6",
    INIT_15 => x"2E2E2E6B7369644D415220676E6974616D726F460D0AB03501E0B70235B03502",
    INIT_16 => x"AAF28E04202164657461636F6C6C6120746F6E206B7369646D6152040D0A0420",
    INIT_17 => x"BD1BDE8E1EDEF7396AF4BDC2F28EF52604C15C0C27018185A65F2ADE8E6AF4BD",
    INIT_18 => x"4C20DEB684A71FDEB646DE8E20DEB701861FDE7FFB265A80A75F4F46DE8E6CF0",
    INIT_19 => x"B70186D7260F8120DEB620DE7C5BF0BD20DEF61FDEB601A70186846C04260F81",
    INIT_1a => x"C6BF86016F846F46DE8E57F0BD0EC6BF8646DE8EC826C0811FDEB61FDE7C20DE",
    INIT_1b => x"03C64F46DE8E5BF0BD0EC64F016F846F46DE8E57F0BD0EC64F46DE8E5BF0BD0E",
    INIT_1c => x"ED204BCC1488ED5349CC1288ED444DCC1088ED4152CC016F846F46DE8E57F0BD",
    INIT_1d => x"01862188ED720ACC2688ED1F88ED0EC6BF861D88ED0101CC1B88ED0100CC1688",
    INIT_1e => x"8646DE8E57F0BD01C64F46DE8E5BF0BD03C64F2588A707862488A707862388A7",
    INIT_1f => x"206C616E7265746E6920676E69746F6F4208085BF07E01C64F01A7558684A7AA",
    INIT_20 => x"26FDD38C81EDA1EC34F48E10E5D38E6AF4BDEDF38E040A0D2E2E2E2E58454C46",
    INIT_21 => x"82F482F4C8DFC2DF82F476F400CD7EF7261EDE8C81EDA1EC4CF48E1000DE8EF7",
    INIT_22 => x"F07E9FF07E6CF07E63F07E5FF07E5BF07E57F07E72F46EF47AF482F47EF482F4",
    INIT_23 => x"9F6E08F89F6E04F89F6E06F89F6E0AF89F6E0CF89F6EC3F07EBFF07EA7F07EA3",
    INIT_24 => x"040A0D2E2E2E2064616F6C7075206B736944204D4F52206C61697265533900F8",
    INIT_25 => x"01C64F1EDEB700866AF4BD83F48E040A0D646564616F4C206B736944204D4F52",
    INIT_26 => x"E0260FC15C20DEF61FDEB626FC17F8265AC0A7EDF4BD5FFEFB1720DEF71FDEB7",
    INIT_27 => x"BD8435E0AB0434068D891F484848480E8D04346AF47EA0F48ED92630814C01C6",
    INIT_28 => x"B7038639018500E0B6390780EB2E1681EF2B11810A2F0981F72B3080FB2928F5",
    INIT_29 => x"DD8D0A2778850826018500E0B629DE7F28DE7F27DEB710863900E0B7118600E0",
    INIT_2a => x"00E0B6023439021A4FDC2627DE7AE12628DE7AE62629DE7A39021C01E0B6E620",
    INIT_2b => x"44204D4F52206D65646F6D580A0D3901E0B70235F120B38DF527788508260285",
    INIT_2c => x"550A0D046574656C706D6F432064616F6C70550A0D0464616F6C7055206B7369",
    INIT_2d => x"B7008625DEBF1AF68E23DEB70186B8FE1772F58E04726F7272452064616F6C70",
    INIT_2e => x"F61FDEB61FFB17F6265AC0A720252B00175FF9FA1720DEF71FDEB701C64F1EDE",
    INIT_2f => x"BE10346DFE169DF58E04FB176AF47E8BF58ED72630814C01C6DE260FC15C20DE",
    INIT_30 => x"F68E06260181903525DEBFED2684ADF1201AF68E4FFF1715860A2823FF1725DE",
    INIT_31 => x"8E062623DEB139FA1C39051A0326188139051A2EFF1706860826048139FA1C3A",
    INIT_32 => x"F68E24DEB7808621DE7FEF2623DEB14339FA1C1AF68E11FF17158639FA1C50F6",
    INIT_33 => x"072621DEB139041AFE1C7BF68E032624DE7A023521DEB721DEBB023439FA1C64",
    INIT_34 => x"4C080839FA1C1AF68EC4FE1715860435031F80C45A301F04340D20068623DE7C",
    INIT_35 => x"46042E4D4F5250206769666E6F63206D6F7266206B736964204D4F522064616F",
    INIT_36 => x"4D4F52040D0A2E2E2E6174616420676E6964616F6C202C434E595320646E756F",
    INIT_37 => x"756F4620746F4E206B736944204D4F52040D0A2E646564616F4C206B73694420",
    INIT_38 => x"00008C1F3015277C8D6C8D00008E20008E105A8D6AF4BD9DF68E040D0A2E646E",
    INIT_39 => x"F71FDEB701C61EDEB74F6AF4BDBFF68E6AF47EF0F68EEB2600008C101F31F326",
    INIT_3a => x"30814C01C6E1260FC15C20DEF61FDEB6ABF917F9265AC0A7678D5F82F91720DE",
    INIT_3b => x"BF46DFBFF92600008C1F3000008EC0E0B70086C0E0B702866AF47EDDF68EDA26",
    INIT_3c => x"FFCC46DF7947DF7948DF793949DF7844C0E0B6C0E0B70086C0E0B701863948DF",
    INIT_3d => x"B2FC17843549DFB6FB265ACE8D08C604343946DFB31055AACC072648DFB31000",
    INIT_3e => x"F4F78EF526F4F78C02300D2780E1E5F78E20C0022F60C1A5FC172086891F7F84",
    INIT_3f => x"000000040D0A3F2054414857ACF55806F750DDF246B2F44C0BF442946E87FC16",

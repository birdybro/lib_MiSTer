    INIT_00 => x"A780A610C6C0DF8E1074FE8E2EFA1AFB1EFB8FFBCEFCB9FC9BFCA1FC61F814F8",
    INIT_01 => x"17431FE4A7D0866AAFDD8C30FB265AE26F0CC65B0117E0DFBF00E08EF9265AA0",
    INIT_02 => x"0317A3FE8E0C0417F62A5A19048B0327856D0DC64FD0DF8E47031784FE8E9F04",
    INIT_03 => x"17408B981F5304175E86092C2081891FF1270D817F84370417B30217AAFE8E2E",
    INIT_04 => x"20F00217ACFE8EF52674FE8C02300F2780E13BFE8E20C0022F60C14704174C04",
    INIT_05 => x"17A4A60F0417A50317211F650217B2FE8E121F2D296B03173B341FBC2094ADC0",
    INIT_06 => x"27A4A1A4A7390F260D8117275E81DD271881E127088111285E0317070417A503",
    INIT_07 => x"0B031705201F30C0DF8E321FA20217BE203F31C2202131E503173F86E8031708",
    INIT_08 => x"279A03170527E4AC011FF0C4201F0634F0C41000C3101F390124E1AC20340629",
    INIT_09 => x"265A8E03172C031780A610C69603172E0317E4AEEE0117B2FE8E103439623203",
    INIT_0a => x"29B70217BC20EE265A7703172E8602237E810425208180A610C6E1AE860317F5",
    INIT_0b => x"3984A73F86A4AFA0A709273F8184A60F271035558DFFFF8E10341A24C0DF8C1E",
    INIT_0c => x"4AAF0427268D1F304AAE431F39FB265A188D08C6E3DF8E104603163F86490317",
    INIT_0d => x"A7A0A7A0A7FF8684A7A4A604263F8184A60A24C0DF8C21AEB9FE16480217068D",
    INIT_0e => x"0186398D46E0B7E086408D393D3139F7265A0427A1ACA0A608C6E3DF8E1039A0",
    INIT_0f => x"178D47E0B7208645E0B744E0B743E0B74F42E0B701862D8D47E0B7EF8641E0B7",

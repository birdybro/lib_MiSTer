    INIT_00 => x"80A608C6023426FF8EC4A6498D1FFF8E292042A6528D1AFF8E2A2046AE5B8D03",
    INIT_01 => x"8D4444444402340235028D023510348235EF265A17FF178200172D860225E468",
    INIT_02 => x"80A64D8D9035048DDFFE8E10340B20028D5C20078B022F3981308B0F84023504",
    INIT_03 => x"86354F0126800017052701C54F0B26618D042702C54FD8F0F6063439F8260481",
    INIT_04 => x"022066001705276200170A2701C510204C00170527478D092702C5D8F0F60434",
    INIT_05 => x"BE84357D0017032701C5358D022702C5D7F0F60434D58DD727D2F07D8435E020",
    INIT_06 => x"F0BE103482350185D0F09FA6023439D2F0B7FF86016D84A7118684A70386D0F0",
    INIT_07 => x"20E0B6023439943501A7FA2702C584E6D0F0BE1434903501A6FA27018584A6D0",
    INIT_08 => x"00CC30E08E943501A7FA2702C584E620E08E14343921E0B6FC27F58D82350185",
    INIT_09 => x"7D30E08E16345986028D1B86D6F07F01E702C6D5F0FD04E703E702A7D3F0FD00",
    INIT_0a => x"101B814100271008819635C5001784A70520098D042420810D20748D0427D6F0",
    INIT_0b => x"0027100B812C0027100C81990027100D814500271016818E0027101A816C0027",
    INIT_0c => x"F0B67400165A3C0027105DD3F0FC9900168300261019C15CD3F0FC51260A8111",
    INIT_0d => x"273DC1D6F0F65800160000CC5B00162500271050814CD3F0B66800164A3327D3",
    INIT_0e => x"39D5F0B70426D5F07D39D6F07F39D6F0B704263D81312754816E002710598116",
    INIT_0f => x"C6D3F0B6168D0000CC1B20E12218C120C0D5F07FD5F0F6ED224F812080D6F07F",

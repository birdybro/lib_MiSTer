    INIT_00 => x"8AE28AE28AE28AE28AE28AE28AE2C1E4C5E4D0E405E5D7E403E5E8E479E038E0",
    INIT_01 => x"C6C07F8E108CE58EC07FCE108AE28AE28AE28AE23EE52FE525E512E58AE28AE2",
    INIT_02 => x"A7D0866AAFDD8C30FB265AE26F0CC6760117D67FBF08808EF9265AA0A780A612",
    INIT_03 => x"17420417BAE58E5704179EE58EC50117A20417DA7FB70386D97FB70386431FE4",
    INIT_04 => x"4DE58E1803176B0417408B981F7204175E86092C2081891FF1270D817F846604",
    INIT_05 => x"E58E121F2D29BA0217C22094ADC6201F0417BCE58EF5268CE58C02300F2780E1",
    INIT_06 => x"271881E12708811128AD0217E10217DA0317A4A6E90217DA0317211FFD0317C2",
    INIT_07 => x"BE203F31C22021310D04173F86C202170827A4A1A4A7390F260D8117275E81DD",
    INIT_08 => x"34F0C41000C3101F390124E1AC203406295B021705201F30C07F8E321F350317",
    INIT_09 => x"630317E4AE860317C2E58E10343962320327A903170527E4AC011FF0C4201F06",
    INIT_0a => x"237E810425208180A610C6E1AE600217F5265A68021761031780A610C6700217",
    INIT_0b => x"C8930317072653817003175F3B341F390128720217BC20EE265A9F03172E8602",
    INIT_0c => x"8C1F29D7011739DA7FF7F22002C8800317072653815D03175F39D97FF7F22002",
    INIT_0d => x"173984A73F86A4AFA0A709273F8184A60F271035DF0017FFFF8E10341B24C07F",
    INIT_0e => x"29950117D901171C2909021739FA265AA1001708C6DB7F8E103E03163F86F301",
    INIT_0f => x"0480B60580B73686431F392020450017CC7FBFF6E18ED27FBFCC7FBED47FBF14",
    INIT_10 => x"80B736860480B70D86341FD47FBF1F301F27D47FBE24273F8184A64AAE170217",
    INIT_11 => x"B73A860580B7328641FE16CC7FBFD27FBE3B0580B73F860780B736860480B605",
    INIT_12 => x"272C8D1F304AAE431F390780B73E860580B736860680B700860480B7FF860780",
    INIT_13 => x"A4A604263F8184A60A24C07F8C21AE08FE16D47FBF00008EB201170C8D4AAF04",
    INIT_14 => x"1186393D3139F7265A0427A1ACA0A608C6DB7F8E1039A0A7A0A7A0A7FF8684A7",
    INIT_15 => x"001726290234CA0017F12631813C2739814F0217F9265381560217D87F7F528D",
    INIT_16 => x"0527E46AE0EB02340C290435B000170434E46AE46AE4EBE0EBE0E610342129B3",
    INIT_17 => x"AC4A2930346F8DE26F0E02161386D87F73058D3F86B327FFC102355FEB2080A7",
    INIT_18 => x"1703E68E64E720C6022320008310062762A3E4ECF901171286E4AF0130462562",
    INIT_19 => x"981F53F526646A72011780A684EB63EB62EB75011762AE820117981F03CB9F01",
    INIT_1a => x"A0A60929188D5D8D3E8610341529188D3965326A8D1486C326E4AC62AF680117",
    INIT_1b => x"10343229088D011F38290E8D438D2D86121F4229088D391035F726E4AC1080A7",
    INIT_1c => x"39811225308164011739E0AB04341E29078D891F484848482829118D903561A7",
    INIT_1d => x"8DF68D8500174B01162086008D39021A39378003224681072541813930800322",
    INIT_1e => x"7E8D3943A70229AB8DDE8D8000173941A70229B78DEA8D8300173944AF0229B3",
    INIT_1f => x"3946AF022979FF17BD8D7A8D3948AF0229858DC88D7C8D394AAF0229908DD38D",
    INIT_20 => x"A10017C2E58E39C4A7808A042971FF17A58D748D3942A702297DFF17B18D778D",
    INIT_21 => x"311F920017C6E58E4A20438D3C8D358D910017C2E58E348D2D8D268D1E8D168D",
    INIT_22 => x"E58E4D2043A6768DE4E58E562041A67F8DEAE58E572044AE880017DEE58E6120",
    INIT_23 => x"42A6528DEFE58E2A2046AE5B8DD8E58E332048AE648DD2E58E3C204AAE6D8DCC",
    INIT_24 => x"265A17FF176A00172D860225E46880A608C60234FBE58EC4A6498DF4E58E2920",
    INIT_25 => x"20078B022F3981308B0F840235048D4444444402340235028D023510348235EF",
    INIT_26 => x"2702C54FDA7FF6063439F826048180A6358D9035048DB4E58E10340B20028D44",
    INIT_27 => x"7F7D8435EE2002203700170527328D092702C5DA7FF6043486354F0126428D04",
    INIT_28 => x"86016D84A7118684A70386D67FBE84352E8D022702C5D97FF60434E38DE527D8",
    INIT_29 => x"1434903501A6FA27018584A6D67FBE103482350185D67F9FA6023439D87FB7FF",
    INIT_2a => x"18E9E315DEE310D2E3040CE40300E402C6E301943501A7FA2702C584E6D67FBE",
    INIT_2b => x"1AE452F7E25074E14FB7E04D9EE24C87E1496BE1470CE1459AE142F4E319BAE3",
    INIT_2c => x"0000FFFFFFFF34E057E273E173E173E173E173E150E35AC7E158D4E15400E153",
    INIT_2d => x"54414857043E040000000A0D04312E31562067754265636172540000000A0D00",
    INIT_2e => x"2020043D59492020043D50552020043D43502020043D5053202004202D20043F",
    INIT_2f => x"4E4948464504203A43432020043D422020043D412020043D50442020043D5849",
    INIT_30 => x"431FCC7F9F6ECA7F9F6EC87F9F6EC67F9F6EC47F9F6EC07F9F6E04315343565A",
    INIT_31 => x"F16E44AEC4EC10340822D07FBC8B300F27FFFF8CCE7FBE49584F4AAF80E64AAE",
    INIT_32 => x"000000000000000000000000000000000000000000000000C27F9F6E42EE1F37",
    INIT_33 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_34 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_35 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_36 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_37 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_38 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_39 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3a => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3b => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3c => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3d => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3e => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_3f => x"0000000000000000000000000000000000000000000000000000000000000000",
